module top_module (
    input [3:0] in,
    output reg [1:0] pos  );

endmodule
